module core_tb();
endmodule