module alu(
    input [31:0] a,
    input [31:0] b,
    input [???:0] func,
    output r,
    output [???:0] flag
);
endmodule