`timescale 1ns/1ns
module queue_tb();
endmodule